/*		 _   / '_/ 
 *		/ ()/)/ /                   
 *                           
 *   design 	:  approximate FP multiplication (binary16 alt & binary8 
 *				   A Transprecision Floating-Point Platform for Ultra-Low Power Computing 
 *				   https://arxiv.org/abs/1711.10374)                 
 *   date		:  21.02.2018                      
 *   version	:  1.0                      
 *                           
 */

