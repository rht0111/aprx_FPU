/*		 _   / '_/ 
 *		/ ()/)/ /                   
 *                           
 *   design 	:  approximate FPU (binary16 alt & binary8 
 *				   A Transprecision Floating-Point Platform for Ultra-Low Power Computing 
 *				   https://arxiv.org/abs/1711.10374
 * 				   https://github.com/pulp-platform/riscv )                 
 *   date		:  21.02.2018                      
 *   version	:  1.0                      
 *                           
 */

